library ieee;
use ieee.std_logic_1164.all;

entity inc_dec_7bits is
    port(
        d_in    : in std_logic_vector(6 downto 0);
        sel     : in std_logic;
        d_out   : out std_logic;
    );
end inc_dec_7bits;

architecture structural of inc_dec_7bits is
    
    
    
    
    begin
    


end structural;